`define INSTRUCT_MEM_SIZE		256
//`define BENCHMARK "../sim/test1_assembly.txt"
//`define BENCHMARK "../sim/CPU_Testbench/test2_alu_assembly.txt"
//`define BENCHMARK "../sim/CPU_Testbench/test3_mem_assembly.txt"
//`define BENCHMARK "../sim/CPU_Testbench/test4_br_assembly.txt"

`timescale 1ns/10ps

module instructmem (
    input	logic	[31:0]	address,
    output	logic	[31:0]	instruction,
    output  logic   instrMemRdy,
    input	logic	clk	// Memory is combinational, but used for error-checking
    );

    assign instrMemRdy = 1'b1;
   
    // Make sure size is a power of two and reasonable.
    initial assert((`INSTRUCT_MEM_SIZE & (`INSTRUCT_MEM_SIZE-1)) == 0 && `INSTRUCT_MEM_SIZE > 4);
    
    // Make sure accesses are reasonable.
    always_ff @(posedge clk) begin
        if (address !== 'x) begin // address or size could be all X's at startup, so ignore this case.
            assert(address[1:0] == 0);	// Makes sure address is aligned.
            assert(address + 3 < `INSTRUCT_MEM_SIZE);	// Make sure address in bounds.
        end
    end
    
    // The data storage itself.
    logic [31:0] mem [`INSTRUCT_MEM_SIZE/4-1:0];
    
    // Load the program - change the filename to pick a different program.
    initial begin
        $readmemb(`BENCHMARK, mem);
        $display("Running benchmark: ", `BENCHMARK);
    end
    
    // Handle the reads.
    integer i;
    always_comb begin
        if (address + 3 >= `INSTRUCT_MEM_SIZE)
            instruction = 'x;
        else
            instruction = mem[address/4];
    end
        
endmodule

module instructmem_testbench ();

    parameter ClockDelay = 5000;

    logic		[63:0]	address;
    logic					clk;
    logic		[31:0]	instruction;
    
    instructmem dut (.address, .instruction, .clk);
    
    initial begin // Set up the clock
        clk <= 0;
        forever #(ClockDelay/2) clk <= ~clk;
    end
    
    integer i;
    initial begin
        // Read every location, including just past the end of the memory.
        for (i=0; i <= `INSTRUCT_MEM_SIZE; i = i + 4) begin
            address <= i;
            @(posedge clk); 
        end
        $stop;
        
    end
endmodule
