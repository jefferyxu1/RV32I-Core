//Adapted from this source: https://download.csdn.net/download/mytlyan/10909630?ops_request_misc=%257B%2522request%255Fid%2522%253A%2522164764800516780269838964%2522%252C%2522scm%2522%253A%252220140713.130102334..%2522%257D&request_id=164764800516780269838964&biz_id=1&utm_medium=distribute.pc_search_result.none-task-download-2~all~sobaiduend~default-2-10909630.142^v2^pc_search_result_control_group,143^v4^register&utm_term=kogge-stone+%E6%A0%91%E5%BD%A2%E5%8A%A0%E6%B3%95%E5%99%A8&spm=1018.2226.3001.4187.3

`timescale 1ns/10ps


`default_nettype none

module dot_operation(p,g,p_1,g_1,p_2,g_2);
    output wire p, g;
    input wire p_1, g_1, p_2, g_2;
    assign p=p_1&p_2;
    assign g=g_2|(p_2&g_1);
endmodule

module get_pg(p,g,a,b);
    output wire p, g;
    input wire a, b;
    assign p=a^b;
    assign g=a&b;
endmodule

// top kogge stone adder top level module
module ksa_top(
    input wire [31:0] a, b,
    input wire cin,     // cin = 0 is addition, cin = 1 is subtraction
    output wire carryOut, overflow, zero, neg,
    output wire [31:0] sum);

    wire [31:0] input_a, input_b;
    assign input_a = a;

    assign input_b = cin ? ~b : b;

    wire c_out_0;
    wire c_out_1;
    wire c_out_2;
    wire c_out_3;
    wire c_out_4;
    wire c_out_5;
    wire c_out_6;
    wire c_out_7;
    wire c_out_8;
    wire c_out_9;
    wire c_out_10;
    wire c_out_11;
    wire c_out_12;
    wire c_out_13;
    wire c_out_14;
    wire c_out_15;
    wire c_out_16;
    wire c_out_17;
    wire c_out_18;
    wire c_out_19;
    wire c_out_20;
    wire c_out_21;
    wire c_out_22;
    wire c_out_23;
    wire c_out_24;
    wire c_out_25;
    wire c_out_26;
    wire c_out_27;
    wire c_out_28;
    wire c_out_29;
    wire c_out_30;
    wire c_out_31;
    wire p_0_0;
    wire g_0_0;
    wire p_1_1;
    wire g_1_1;
    wire p_2_2;
    wire g_2_2;
    wire p_3_3;
    wire g_3_3;
    wire p_4_4;
    wire g_4_4;
    wire p_5_5;
    wire g_5_5;
    wire p_6_6;
    wire g_6_6;
    wire p_7_7;
    wire g_7_7;
    wire p_8_8;
    wire g_8_8;
    wire p_9_9;
    wire g_9_9;
    wire p_10_10;
    wire g_10_10;
    wire p_11_11;
    wire g_11_11;
    wire p_12_12;
    wire g_12_12;
    wire p_13_13;
    wire g_13_13;
    wire p_14_14;
    wire g_14_14;
    wire p_15_15;
    wire g_15_15;
    wire p_16_16;
    wire g_16_16;
    wire p_17_17;
    wire g_17_17;
    wire p_18_18;
    wire g_18_18;
    wire p_19_19;
    wire g_19_19;
    wire p_20_20;
    wire g_20_20;
    wire p_21_21;
    wire g_21_21;
    wire p_22_22;
    wire g_22_22;
    wire p_23_23;
    wire g_23_23;
    wire p_24_24;
    wire g_24_24;
    wire p_25_25;
    wire g_25_25;
    wire p_26_26;
    wire g_26_26;
    wire p_27_27;
    wire g_27_27;
    wire p_28_28;
    wire g_28_28;
    wire p_29_29;
    wire g_29_29;
    wire p_30_30;
    wire g_30_30;
    wire p_31_31;
    wire g_31_31;
//get pg

    get_pg get_0_0(.p(p_0_0),.g(g_0_0),.a(input_a[0]),.b(input_b[0]));
    get_pg get_1_1(.p(p_1_1),.g(g_1_1),.a(input_a[1]),.b(input_b[1]));
    get_pg get_2_2(.p(p_2_2),.g(g_2_2),.a(input_a[2]),.b(input_b[2]));
    get_pg get_3_3(.p(p_3_3),.g(g_3_3),.a(input_a[3]),.b(input_b[3]));
    get_pg get_4_4(.p(p_4_4),.g(g_4_4),.a(input_a[4]),.b(input_b[4]));
    get_pg get_5_5(.p(p_5_5),.g(g_5_5),.a(input_a[5]),.b(input_b[5]));
    get_pg get_6_6(.p(p_6_6),.g(g_6_6),.a(input_a[6]),.b(input_b[6]));
    get_pg get_7_7(.p(p_7_7),.g(g_7_7),.a(input_a[7]),.b(input_b[7]));
    get_pg get_8_8(.p(p_8_8),.g(g_8_8),.a(input_a[8]),.b(input_b[8]));
    get_pg get_9_9(.p(p_9_9),.g(g_9_9),.a(input_a[9]),.b(input_b[9]));
    get_pg get_10_10(.p(p_10_10),.g(g_10_10),.a(input_a[10]),.b(input_b[10]));
    get_pg get_11_11(.p(p_11_11),.g(g_11_11),.a(input_a[11]),.b(input_b[11]));
    get_pg get_12_12(.p(p_12_12),.g(g_12_12),.a(input_a[12]),.b(input_b[12]));
    get_pg get_13_13(.p(p_13_13),.g(g_13_13),.a(input_a[13]),.b(input_b[13]));
    get_pg get_14_14(.p(p_14_14),.g(g_14_14),.a(input_a[14]),.b(input_b[14]));
    get_pg get_15_15(.p(p_15_15),.g(g_15_15),.a(input_a[15]),.b(input_b[15]));
    get_pg get_16_16(.p(p_16_16),.g(g_16_16),.a(input_a[16]),.b(input_b[16]));
    get_pg get_17_17(.p(p_17_17),.g(g_17_17),.a(input_a[17]),.b(input_b[17]));
    get_pg get_18_18(.p(p_18_18),.g(g_18_18),.a(input_a[18]),.b(input_b[18]));
    get_pg get_19_19(.p(p_19_19),.g(g_19_19),.a(input_a[19]),.b(input_b[19]));
    get_pg get_20_20(.p(p_20_20),.g(g_20_20),.a(input_a[20]),.b(input_b[20]));
    get_pg get_21_21(.p(p_21_21),.g(g_21_21),.a(input_a[21]),.b(input_b[21]));
    get_pg get_22_22(.p(p_22_22),.g(g_22_22),.a(input_a[22]),.b(input_b[22]));
    get_pg get_23_23(.p(p_23_23),.g(g_23_23),.a(input_a[23]),.b(input_b[23]));
    get_pg get_24_24(.p(p_24_24),.g(g_24_24),.a(input_a[24]),.b(input_b[24]));
    get_pg get_25_25(.p(p_25_25),.g(g_25_25),.a(input_a[25]),.b(input_b[25]));
    get_pg get_26_26(.p(p_26_26),.g(g_26_26),.a(input_a[26]),.b(input_b[26]));
    get_pg get_27_27(.p(p_27_27),.g(g_27_27),.a(input_a[27]),.b(input_b[27]));
    get_pg get_28_28(.p(p_28_28),.g(g_28_28),.a(input_a[28]),.b(input_b[28]));
    get_pg get_29_29(.p(p_29_29),.g(g_29_29),.a(input_a[29]),.b(input_b[29]));
    get_pg get_30_30(.p(p_30_30),.g(g_30_30),.a(input_a[30]),.b(input_b[30]));
    get_pg get_31_31(.p(p_31_31),.g(g_31_31),.a(input_a[31]),.b(input_b[31]));


    wire p_0_1;
    wire g_0_1;
    dot_operation get_0_1(.p(p_0_1),.g(g_0_1),.p_1(p_0_0),.g_1(g_0_0),.p_2(p_1_1),.g_2(g_1_1));
    wire p_1_2;
    wire g_1_2;
    dot_operation get_1_2(.p(p_1_2),.g(g_1_2),.p_1(p_1_1),.g_1(g_1_1),.p_2(p_2_2),.g_2(g_2_2));
    wire p_2_3;
    wire g_2_3;
    dot_operation get_2_3(.p(p_2_3),.g(g_2_3),.p_1(p_2_2),.g_1(g_2_2),.p_2(p_3_3),.g_2(g_3_3));
    wire p_3_4;
    wire g_3_4;
    dot_operation get_3_4(.p(p_3_4),.g(g_3_4),.p_1(p_3_3),.g_1(g_3_3),.p_2(p_4_4),.g_2(g_4_4));
    wire p_4_5;
    wire g_4_5;
    dot_operation get_4_5(.p(p_4_5),.g(g_4_5),.p_1(p_4_4),.g_1(g_4_4),.p_2(p_5_5),.g_2(g_5_5));
    wire p_5_6;
    wire g_5_6;
    dot_operation get_5_6(.p(p_5_6),.g(g_5_6),.p_1(p_5_5),.g_1(g_5_5),.p_2(p_6_6),.g_2(g_6_6));
    wire p_6_7;
    wire g_6_7;
    dot_operation get_6_7(.p(p_6_7),.g(g_6_7),.p_1(p_6_6),.g_1(g_6_6),.p_2(p_7_7),.g_2(g_7_7));
    wire p_7_8;
    wire g_7_8;
    dot_operation get_7_8(.p(p_7_8),.g(g_7_8),.p_1(p_7_7),.g_1(g_7_7),.p_2(p_8_8),.g_2(g_8_8));
    wire p_8_9;
    wire g_8_9;
    dot_operation get_8_9(.p(p_8_9),.g(g_8_9),.p_1(p_8_8),.g_1(g_8_8),.p_2(p_9_9),.g_2(g_9_9));
    wire p_9_10;
    wire g_9_10;
    dot_operation get_9_10(.p(p_9_10),.g(g_9_10),.p_1(p_9_9),.g_1(g_9_9),.p_2(p_10_10),.g_2(g_10_10));
    wire p_10_11;
    wire g_10_11;
    dot_operation get_10_11(.p(p_10_11),.g(g_10_11),.p_1(p_10_10),.g_1(g_10_10),.p_2(p_11_11),.g_2(g_11_11));
    wire p_11_12;
    wire g_11_12;
    dot_operation get_11_12(.p(p_11_12),.g(g_11_12),.p_1(p_11_11),.g_1(g_11_11),.p_2(p_12_12),.g_2(g_12_12));
    wire p_12_13;
    wire g_12_13;
    dot_operation get_12_13(.p(p_12_13),.g(g_12_13),.p_1(p_12_12),.g_1(g_12_12),.p_2(p_13_13),.g_2(g_13_13));
    wire p_13_14;
    wire g_13_14;
    dot_operation get_13_14(.p(p_13_14),.g(g_13_14),.p_1(p_13_13),.g_1(g_13_13),.p_2(p_14_14),.g_2(g_14_14));
    wire p_14_15;
    wire g_14_15;
    dot_operation get_14_15(.p(p_14_15),.g(g_14_15),.p_1(p_14_14),.g_1(g_14_14),.p_2(p_15_15),.g_2(g_15_15));
    wire p_15_16;
    wire g_15_16;
    dot_operation get_15_16(.p(p_15_16),.g(g_15_16),.p_1(p_15_15),.g_1(g_15_15),.p_2(p_16_16),.g_2(g_16_16));
    wire p_16_17;
    wire g_16_17;
    dot_operation get_16_17(.p(p_16_17),.g(g_16_17),.p_1(p_16_16),.g_1(g_16_16),.p_2(p_17_17),.g_2(g_17_17));
    wire p_17_18;
    wire g_17_18;
    dot_operation get_17_18(.p(p_17_18),.g(g_17_18),.p_1(p_17_17),.g_1(g_17_17),.p_2(p_18_18),.g_2(g_18_18));
    wire p_18_19;
    wire g_18_19;
    dot_operation get_18_19(.p(p_18_19),.g(g_18_19),.p_1(p_18_18),.g_1(g_18_18),.p_2(p_19_19),.g_2(g_19_19));
    wire p_19_20;
    wire g_19_20;
    dot_operation get_19_20(.p(p_19_20),.g(g_19_20),.p_1(p_19_19),.g_1(g_19_19),.p_2(p_20_20),.g_2(g_20_20));
    wire p_20_21;
    wire g_20_21;
    dot_operation get_20_21(.p(p_20_21),.g(g_20_21),.p_1(p_20_20),.g_1(g_20_20),.p_2(p_21_21),.g_2(g_21_21));
    wire p_21_22;
    wire g_21_22;
    dot_operation get_21_22(.p(p_21_22),.g(g_21_22),.p_1(p_21_21),.g_1(g_21_21),.p_2(p_22_22),.g_2(g_22_22));
    wire p_22_23;
    wire g_22_23;
    dot_operation get_22_23(.p(p_22_23),.g(g_22_23),.p_1(p_22_22),.g_1(g_22_22),.p_2(p_23_23),.g_2(g_23_23));
    wire p_23_24;
    wire g_23_24;
    dot_operation get_23_24(.p(p_23_24),.g(g_23_24),.p_1(p_23_23),.g_1(g_23_23),.p_2(p_24_24),.g_2(g_24_24));
    wire p_24_25;
    wire g_24_25;
    dot_operation get_24_25(.p(p_24_25),.g(g_24_25),.p_1(p_24_24),.g_1(g_24_24),.p_2(p_25_25),.g_2(g_25_25));
    wire p_25_26;
    wire g_25_26;
    dot_operation get_25_26(.p(p_25_26),.g(g_25_26),.p_1(p_25_25),.g_1(g_25_25),.p_2(p_26_26),.g_2(g_26_26));
    wire p_26_27;
    wire g_26_27;
    dot_operation get_26_27(.p(p_26_27),.g(g_26_27),.p_1(p_26_26),.g_1(g_26_26),.p_2(p_27_27),.g_2(g_27_27));
    wire p_27_28;
    wire g_27_28;
    dot_operation get_27_28(.p(p_27_28),.g(g_27_28),.p_1(p_27_27),.g_1(g_27_27),.p_2(p_28_28),.g_2(g_28_28));
    wire p_28_29;
    wire g_28_29;
    dot_operation get_28_29(.p(p_28_29),.g(g_28_29),.p_1(p_28_28),.g_1(g_28_28),.p_2(p_29_29),.g_2(g_29_29));
    wire p_29_30;
    wire g_29_30;
    dot_operation get_29_30(.p(p_29_30),.g(g_29_30),.p_1(p_29_29),.g_1(g_29_29),.p_2(p_30_30),.g_2(g_30_30));
    wire p_30_31;
    wire g_30_31;
    dot_operation get_30_31(.p(p_30_31),.g(g_30_31),.p_1(p_30_30),.g_1(g_30_30),.p_2(p_31_31),.g_2(g_31_31));
    wire p_0_2;
    wire g_0_2;
    dot_operation get_0_2(.p(p_0_2),.g(g_0_2),.p_1(p_0_0),.g_1(g_0_0),.p_2(p_1_2),.g_2(g_1_2));
    wire p_0_3;
    wire g_0_3;
    dot_operation get_0_3(.p(p_0_3),.g(g_0_3),.p_1(p_0_1),.g_1(g_0_1),.p_2(p_2_3),.g_2(g_2_3));
    wire p_1_4;
    wire g_1_4;
    dot_operation get_1_4(.p(p_1_4),.g(g_1_4),.p_1(p_1_2),.g_1(g_1_2),.p_2(p_3_4),.g_2(g_3_4));
    wire p_2_5;
    wire g_2_5;
    dot_operation get_2_5(.p(p_2_5),.g(g_2_5),.p_1(p_2_3),.g_1(g_2_3),.p_2(p_4_5),.g_2(g_4_5));
    wire p_3_6;
    wire g_3_6;
    dot_operation get_3_6(.p(p_3_6),.g(g_3_6),.p_1(p_3_4),.g_1(g_3_4),.p_2(p_5_6),.g_2(g_5_6));
    wire p_4_7;
    wire g_4_7;
    dot_operation get_4_7(.p(p_4_7),.g(g_4_7),.p_1(p_4_5),.g_1(g_4_5),.p_2(p_6_7),.g_2(g_6_7));
    wire p_5_8;
    wire g_5_8;
    dot_operation get_5_8(.p(p_5_8),.g(g_5_8),.p_1(p_5_6),.g_1(g_5_6),.p_2(p_7_8),.g_2(g_7_8));
    wire p_6_9;
    wire g_6_9;
    dot_operation get_6_9(.p(p_6_9),.g(g_6_9),.p_1(p_6_7),.g_1(g_6_7),.p_2(p_8_9),.g_2(g_8_9));
    wire p_7_10;
    wire g_7_10;
    dot_operation get_7_10(.p(p_7_10),.g(g_7_10),.p_1(p_7_8),.g_1(g_7_8),.p_2(p_9_10),.g_2(g_9_10));
    wire p_8_11;
    wire g_8_11;
    dot_operation get_8_11(.p(p_8_11),.g(g_8_11),.p_1(p_8_9),.g_1(g_8_9),.p_2(p_10_11),.g_2(g_10_11));
    wire p_9_12;
    wire g_9_12;
    dot_operation get_9_12(.p(p_9_12),.g(g_9_12),.p_1(p_9_10),.g_1(g_9_10),.p_2(p_11_12),.g_2(g_11_12));
    wire p_10_13;
    wire g_10_13;
    dot_operation get_10_13(.p(p_10_13),.g(g_10_13),.p_1(p_10_11),.g_1(g_10_11),.p_2(p_12_13),.g_2(g_12_13));
    wire p_11_14;
    wire g_11_14;
    dot_operation get_11_14(.p(p_11_14),.g(g_11_14),.p_1(p_11_12),.g_1(g_11_12),.p_2(p_13_14),.g_2(g_13_14));
    wire p_12_15;
    wire g_12_15;
    dot_operation get_12_15(.p(p_12_15),.g(g_12_15),.p_1(p_12_13),.g_1(g_12_13),.p_2(p_14_15),.g_2(g_14_15));
    wire p_13_16;
    wire g_13_16;
    dot_operation get_13_16(.p(p_13_16),.g(g_13_16),.p_1(p_13_14),.g_1(g_13_14),.p_2(p_15_16),.g_2(g_15_16));
    wire p_14_17;
    wire g_14_17;
    dot_operation get_14_17(.p(p_14_17),.g(g_14_17),.p_1(p_14_15),.g_1(g_14_15),.p_2(p_16_17),.g_2(g_16_17));
    wire p_15_18;
    wire g_15_18;
    dot_operation get_15_18(.p(p_15_18),.g(g_15_18),.p_1(p_15_16),.g_1(g_15_16),.p_2(p_17_18),.g_2(g_17_18));
    wire p_16_19;
    wire g_16_19;
    dot_operation get_16_19(.p(p_16_19),.g(g_16_19),.p_1(p_16_17),.g_1(g_16_17),.p_2(p_18_19),.g_2(g_18_19));
    wire p_17_20;
    wire g_17_20;
    dot_operation get_17_20(.p(p_17_20),.g(g_17_20),.p_1(p_17_18),.g_1(g_17_18),.p_2(p_19_20),.g_2(g_19_20));
    wire p_18_21;
    wire g_18_21;
    dot_operation get_18_21(.p(p_18_21),.g(g_18_21),.p_1(p_18_19),.g_1(g_18_19),.p_2(p_20_21),.g_2(g_20_21));
    wire p_19_22;
    wire g_19_22;
    dot_operation get_19_22(.p(p_19_22),.g(g_19_22),.p_1(p_19_20),.g_1(g_19_20),.p_2(p_21_22),.g_2(g_21_22));
    wire p_20_23;
    wire g_20_23;
    dot_operation get_20_23(.p(p_20_23),.g(g_20_23),.p_1(p_20_21),.g_1(g_20_21),.p_2(p_22_23),.g_2(g_22_23));
    wire p_21_24;
    wire g_21_24;
    dot_operation get_21_24(.p(p_21_24),.g(g_21_24),.p_1(p_21_22),.g_1(g_21_22),.p_2(p_23_24),.g_2(g_23_24));
    wire p_22_25;
    wire g_22_25;
    dot_operation get_22_25(.p(p_22_25),.g(g_22_25),.p_1(p_22_23),.g_1(g_22_23),.p_2(p_24_25),.g_2(g_24_25));
    wire p_23_26;
    wire g_23_26;
    dot_operation get_23_26(.p(p_23_26),.g(g_23_26),.p_1(p_23_24),.g_1(g_23_24),.p_2(p_25_26),.g_2(g_25_26));
    wire p_24_27;
    wire g_24_27;
    dot_operation get_24_27(.p(p_24_27),.g(g_24_27),.p_1(p_24_25),.g_1(g_24_25),.p_2(p_26_27),.g_2(g_26_27));
    wire p_25_28;
    wire g_25_28;
    dot_operation get_25_28(.p(p_25_28),.g(g_25_28),.p_1(p_25_26),.g_1(g_25_26),.p_2(p_27_28),.g_2(g_27_28));
    wire p_26_29;
    wire g_26_29;
    dot_operation get_26_29(.p(p_26_29),.g(g_26_29),.p_1(p_26_27),.g_1(g_26_27),.p_2(p_28_29),.g_2(g_28_29));
    wire p_27_30;
    wire g_27_30;
    dot_operation get_27_30(.p(p_27_30),.g(g_27_30),.p_1(p_27_28),.g_1(g_27_28),.p_2(p_29_30),.g_2(g_29_30));
    wire p_28_31;
    wire g_28_31;
    dot_operation get_28_31(.p(p_28_31),.g(g_28_31),.p_1(p_28_29),.g_1(g_28_29),.p_2(p_30_31),.g_2(g_30_31));
    wire p_0_4;
    wire g_0_4;
    dot_operation get_0_4(.p(p_0_4),.g(g_0_4),.p_1(p_0_0),.g_1(g_0_0),.p_2(p_1_4),.g_2(g_1_4));
    wire p_0_5;
    wire g_0_5;
    dot_operation get_0_5(.p(p_0_5),.g(g_0_5),.p_1(p_0_1),.g_1(g_0_1),.p_2(p_2_5),.g_2(g_2_5));
    wire p_0_6;
    wire g_0_6;
    dot_operation get_0_6(.p(p_0_6),.g(g_0_6),.p_1(p_0_2),.g_1(g_0_2),.p_2(p_3_6),.g_2(g_3_6));
    wire p_0_7;
    wire g_0_7;
    dot_operation get_0_7(.p(p_0_7),.g(g_0_7),.p_1(p_0_3),.g_1(g_0_3),.p_2(p_4_7),.g_2(g_4_7));
    wire p_1_8;
    wire g_1_8;
    dot_operation get_1_8(.p(p_1_8),.g(g_1_8),.p_1(p_1_4),.g_1(g_1_4),.p_2(p_5_8),.g_2(g_5_8));
    wire p_2_9;
    wire g_2_9;
    dot_operation get_2_9(.p(p_2_9),.g(g_2_9),.p_1(p_2_5),.g_1(g_2_5),.p_2(p_6_9),.g_2(g_6_9));
    wire p_3_10;
    wire g_3_10;
    dot_operation get_3_10(.p(p_3_10),.g(g_3_10),.p_1(p_3_6),.g_1(g_3_6),.p_2(p_7_10),.g_2(g_7_10));
    wire p_4_11;
    wire g_4_11;
    dot_operation get_4_11(.p(p_4_11),.g(g_4_11),.p_1(p_4_7),.g_1(g_4_7),.p_2(p_8_11),.g_2(g_8_11));
    wire p_5_12;
    wire g_5_12;
    dot_operation get_5_12(.p(p_5_12),.g(g_5_12),.p_1(p_5_8),.g_1(g_5_8),.p_2(p_9_12),.g_2(g_9_12));
    wire p_6_13;
    wire g_6_13;
    dot_operation get_6_13(.p(p_6_13),.g(g_6_13),.p_1(p_6_9),.g_1(g_6_9),.p_2(p_10_13),.g_2(g_10_13));
    wire p_7_14;
    wire g_7_14;
    dot_operation get_7_14(.p(p_7_14),.g(g_7_14),.p_1(p_7_10),.g_1(g_7_10),.p_2(p_11_14),.g_2(g_11_14));
    wire p_8_15;
    wire g_8_15;
    dot_operation get_8_15(.p(p_8_15),.g(g_8_15),.p_1(p_8_11),.g_1(g_8_11),.p_2(p_12_15),.g_2(g_12_15));
    wire p_9_16;
    wire g_9_16;
    dot_operation get_9_16(.p(p_9_16),.g(g_9_16),.p_1(p_9_12),.g_1(g_9_12),.p_2(p_13_16),.g_2(g_13_16));
    wire p_10_17;
    wire g_10_17;
    dot_operation get_10_17(.p(p_10_17),.g(g_10_17),.p_1(p_10_13),.g_1(g_10_13),.p_2(p_14_17),.g_2(g_14_17));
    wire p_11_18;
    wire g_11_18;
    dot_operation get_11_18(.p(p_11_18),.g(g_11_18),.p_1(p_11_14),.g_1(g_11_14),.p_2(p_15_18),.g_2(g_15_18));
    wire p_12_19;
    wire g_12_19;
    dot_operation get_12_19(.p(p_12_19),.g(g_12_19),.p_1(p_12_15),.g_1(g_12_15),.p_2(p_16_19),.g_2(g_16_19));
    wire p_13_20;
    wire g_13_20;
    dot_operation get_13_20(.p(p_13_20),.g(g_13_20),.p_1(p_13_16),.g_1(g_13_16),.p_2(p_17_20),.g_2(g_17_20));
    wire p_14_21;
    wire g_14_21;
    dot_operation get_14_21(.p(p_14_21),.g(g_14_21),.p_1(p_14_17),.g_1(g_14_17),.p_2(p_18_21),.g_2(g_18_21));
    wire p_15_22;
    wire g_15_22;
    dot_operation get_15_22(.p(p_15_22),.g(g_15_22),.p_1(p_15_18),.g_1(g_15_18),.p_2(p_19_22),.g_2(g_19_22));
    wire p_16_23;
    wire g_16_23;
    dot_operation get_16_23(.p(p_16_23),.g(g_16_23),.p_1(p_16_19),.g_1(g_16_19),.p_2(p_20_23),.g_2(g_20_23));
    wire p_17_24;
    wire g_17_24;
    dot_operation get_17_24(.p(p_17_24),.g(g_17_24),.p_1(p_17_20),.g_1(g_17_20),.p_2(p_21_24),.g_2(g_21_24));
    wire p_18_25;
    wire g_18_25;
    dot_operation get_18_25(.p(p_18_25),.g(g_18_25),.p_1(p_18_21),.g_1(g_18_21),.p_2(p_22_25),.g_2(g_22_25));
    wire p_19_26;
    wire g_19_26;
    dot_operation get_19_26(.p(p_19_26),.g(g_19_26),.p_1(p_19_22),.g_1(g_19_22),.p_2(p_23_26),.g_2(g_23_26));
    wire p_20_27;
    wire g_20_27;
    dot_operation get_20_27(.p(p_20_27),.g(g_20_27),.p_1(p_20_23),.g_1(g_20_23),.p_2(p_24_27),.g_2(g_24_27));
    wire p_21_28;
    wire g_21_28;
    dot_operation get_21_28(.p(p_21_28),.g(g_21_28),.p_1(p_21_24),.g_1(g_21_24),.p_2(p_25_28),.g_2(g_25_28));
    wire p_22_29;
    wire g_22_29;
    dot_operation get_22_29(.p(p_22_29),.g(g_22_29),.p_1(p_22_25),.g_1(g_22_25),.p_2(p_26_29),.g_2(g_26_29));
    wire p_23_30;
    wire g_23_30;
    dot_operation get_23_30(.p(p_23_30),.g(g_23_30),.p_1(p_23_26),.g_1(g_23_26),.p_2(p_27_30),.g_2(g_27_30));
    wire p_24_31;
    wire g_24_31;
    dot_operation get_24_31(.p(p_24_31),.g(g_24_31),.p_1(p_24_27),.g_1(g_24_27),.p_2(p_28_31),.g_2(g_28_31));
    wire p_0_8;
    wire g_0_8;
    dot_operation get_0_8(.p(p_0_8),.g(g_0_8),.p_1(p_0_0),.g_1(g_0_0),.p_2(p_1_8),.g_2(g_1_8));
    wire p_0_9;
    wire g_0_9;
    dot_operation get_0_9(.p(p_0_9),.g(g_0_9),.p_1(p_0_1),.g_1(g_0_1),.p_2(p_2_9),.g_2(g_2_9));
    wire p_0_10;
    wire g_0_10;
    dot_operation get_0_10(.p(p_0_10),.g(g_0_10),.p_1(p_0_2),.g_1(g_0_2),.p_2(p_3_10),.g_2(g_3_10));
    wire p_0_11;
    wire g_0_11;
    dot_operation get_0_11(.p(p_0_11),.g(g_0_11),.p_1(p_0_3),.g_1(g_0_3),.p_2(p_4_11),.g_2(g_4_11));
    wire p_0_12;
    wire g_0_12;
    dot_operation get_0_12(.p(p_0_12),.g(g_0_12),.p_1(p_0_4),.g_1(g_0_4),.p_2(p_5_12),.g_2(g_5_12));
    wire p_0_13;
    wire g_0_13;
    dot_operation get_0_13(.p(p_0_13),.g(g_0_13),.p_1(p_0_5),.g_1(g_0_5),.p_2(p_6_13),.g_2(g_6_13));
    wire p_0_14;
    wire g_0_14;
    dot_operation get_0_14(.p(p_0_14),.g(g_0_14),.p_1(p_0_6),.g_1(g_0_6),.p_2(p_7_14),.g_2(g_7_14));
    wire p_0_15;
    wire g_0_15;
    dot_operation get_0_15(.p(p_0_15),.g(g_0_15),.p_1(p_0_7),.g_1(g_0_7),.p_2(p_8_15),.g_2(g_8_15));
    wire p_1_16;
    wire g_1_16;
    dot_operation get_1_16(.p(p_1_16),.g(g_1_16),.p_1(p_1_8),.g_1(g_1_8),.p_2(p_9_16),.g_2(g_9_16));
    wire p_2_17;
    wire g_2_17;
    dot_operation get_2_17(.p(p_2_17),.g(g_2_17),.p_1(p_2_9),.g_1(g_2_9),.p_2(p_10_17),.g_2(g_10_17));
    wire p_3_18;
    wire g_3_18;
    dot_operation get_3_18(.p(p_3_18),.g(g_3_18),.p_1(p_3_10),.g_1(g_3_10),.p_2(p_11_18),.g_2(g_11_18));
    wire p_4_19;
    wire g_4_19;
    dot_operation get_4_19(.p(p_4_19),.g(g_4_19),.p_1(p_4_11),.g_1(g_4_11),.p_2(p_12_19),.g_2(g_12_19));
    wire p_5_20;
    wire g_5_20;
    dot_operation get_5_20(.p(p_5_20),.g(g_5_20),.p_1(p_5_12),.g_1(g_5_12),.p_2(p_13_20),.g_2(g_13_20));
    wire p_6_21;
    wire g_6_21;
    dot_operation get_6_21(.p(p_6_21),.g(g_6_21),.p_1(p_6_13),.g_1(g_6_13),.p_2(p_14_21),.g_2(g_14_21));
    wire p_7_22;
    wire g_7_22;
    dot_operation get_7_22(.p(p_7_22),.g(g_7_22),.p_1(p_7_14),.g_1(g_7_14),.p_2(p_15_22),.g_2(g_15_22));
    wire p_8_23;
    wire g_8_23;
    dot_operation get_8_23(.p(p_8_23),.g(g_8_23),.p_1(p_8_15),.g_1(g_8_15),.p_2(p_16_23),.g_2(g_16_23));
    wire p_9_24;
    wire g_9_24;
    dot_operation get_9_24(.p(p_9_24),.g(g_9_24),.p_1(p_9_16),.g_1(g_9_16),.p_2(p_17_24),.g_2(g_17_24));
    wire p_10_25;
    wire g_10_25;
    dot_operation get_10_25(.p(p_10_25),.g(g_10_25),.p_1(p_10_17),.g_1(g_10_17),.p_2(p_18_25),.g_2(g_18_25));
    wire p_11_26;
    wire g_11_26;
    dot_operation get_11_26(.p(p_11_26),.g(g_11_26),.p_1(p_11_18),.g_1(g_11_18),.p_2(p_19_26),.g_2(g_19_26));
    wire p_12_27;
    wire g_12_27;
    dot_operation get_12_27(.p(p_12_27),.g(g_12_27),.p_1(p_12_19),.g_1(g_12_19),.p_2(p_20_27),.g_2(g_20_27));
    wire p_13_28;
    wire g_13_28;
    dot_operation get_13_28(.p(p_13_28),.g(g_13_28),.p_1(p_13_20),.g_1(g_13_20),.p_2(p_21_28),.g_2(g_21_28));
    wire p_14_29;
    wire g_14_29;
    dot_operation get_14_29(.p(p_14_29),.g(g_14_29),.p_1(p_14_21),.g_1(g_14_21),.p_2(p_22_29),.g_2(g_22_29));
    wire p_15_30;
    wire g_15_30;
    dot_operation get_15_30(.p(p_15_30),.g(g_15_30),.p_1(p_15_22),.g_1(g_15_22),.p_2(p_23_30),.g_2(g_23_30));
    wire p_16_31;
    wire g_16_31;
    dot_operation get_16_31(.p(p_16_31),.g(g_16_31),.p_1(p_16_23),.g_1(g_16_23),.p_2(p_24_31),.g_2(g_24_31));
    wire p_0_16;
    wire g_0_16;
    dot_operation get_0_16(.p(p_0_16),.g(g_0_16),.p_1(p_0_0),.g_1(g_0_0),.p_2(p_1_16),.g_2(g_1_16));
    wire p_0_17;
    wire g_0_17;
    dot_operation get_0_17(.p(p_0_17),.g(g_0_17),.p_1(p_0_1),.g_1(g_0_1),.p_2(p_2_17),.g_2(g_2_17));
    wire p_0_18;
    wire g_0_18;
    dot_operation get_0_18(.p(p_0_18),.g(g_0_18),.p_1(p_0_2),.g_1(g_0_2),.p_2(p_3_18),.g_2(g_3_18));
    wire p_0_19;
    wire g_0_19;
    dot_operation get_0_19(.p(p_0_19),.g(g_0_19),.p_1(p_0_3),.g_1(g_0_3),.p_2(p_4_19),.g_2(g_4_19));
    wire p_0_20;
    wire g_0_20;
    dot_operation get_0_20(.p(p_0_20),.g(g_0_20),.p_1(p_0_4),.g_1(g_0_4),.p_2(p_5_20),.g_2(g_5_20));
    wire p_0_21;
    wire g_0_21;
    dot_operation get_0_21(.p(p_0_21),.g(g_0_21),.p_1(p_0_5),.g_1(g_0_5),.p_2(p_6_21),.g_2(g_6_21));
    wire p_0_22;
    wire g_0_22;
    dot_operation get_0_22(.p(p_0_22),.g(g_0_22),.p_1(p_0_6),.g_1(g_0_6),.p_2(p_7_22),.g_2(g_7_22));
    wire p_0_23;
    wire g_0_23;
    dot_operation get_0_23(.p(p_0_23),.g(g_0_23),.p_1(p_0_7),.g_1(g_0_7),.p_2(p_8_23),.g_2(g_8_23));
    wire p_0_24;
    wire g_0_24;
    dot_operation get_0_24(.p(p_0_24),.g(g_0_24),.p_1(p_0_8),.g_1(g_0_8),.p_2(p_9_24),.g_2(g_9_24));
    wire p_0_25;
    wire g_0_25;
    dot_operation get_0_25(.p(p_0_25),.g(g_0_25),.p_1(p_0_9),.g_1(g_0_9),.p_2(p_10_25),.g_2(g_10_25));
    wire p_0_26;
    wire g_0_26;
    dot_operation get_0_26(.p(p_0_26),.g(g_0_26),.p_1(p_0_10),.g_1(g_0_10),.p_2(p_11_26),.g_2(g_11_26));
    wire p_0_27;
    wire g_0_27;
    dot_operation get_0_27(.p(p_0_27),.g(g_0_27),.p_1(p_0_11),.g_1(g_0_11),.p_2(p_12_27),.g_2(g_12_27));
    wire p_0_28;
    wire g_0_28;
    dot_operation get_0_28(.p(p_0_28),.g(g_0_28),.p_1(p_0_12),.g_1(g_0_12),.p_2(p_13_28),.g_2(g_13_28));
    wire p_0_29;
    wire g_0_29;
    dot_operation get_0_29(.p(p_0_29),.g(g_0_29),.p_1(p_0_13),.g_1(g_0_13),.p_2(p_14_29),.g_2(g_14_29));
    wire p_0_30;
    wire g_0_30;
    dot_operation get_0_30(.p(p_0_30),.g(g_0_30),.p_1(p_0_14),.g_1(g_0_14),.p_2(p_15_30),.g_2(g_15_30));
    wire p_0_31;
    wire g_0_31;
    dot_operation get_0_31(.p(p_0_31),.g(g_0_31),.p_1(p_0_15),.g_1(g_0_15),.p_2(p_16_31),.g_2(g_16_31));
    assign c_out_0=g_0_0|(p_0_0&cin);
    assign c_out_1=g_0_1|(p_0_1&cin);
    assign c_out_2=g_0_2|(p_0_2&cin);
    assign c_out_3=g_0_3|(p_0_3&cin);
    assign c_out_4=g_0_4|(p_0_4&cin);
    assign c_out_5=g_0_5|(p_0_5&cin);
    assign c_out_6=g_0_6|(p_0_6&cin);
    assign c_out_7=g_0_7|(p_0_7&cin);
    assign c_out_8=g_0_8|(p_0_8&cin);
    assign c_out_9=g_0_9|(p_0_9&cin);
    assign c_out_10=g_0_10|(p_0_10&cin);
    assign c_out_11=g_0_11|(p_0_11&cin);
    assign c_out_12=g_0_12|(p_0_12&cin);
    assign c_out_13=g_0_13|(p_0_13&cin);
    assign c_out_14=g_0_14|(p_0_14&cin);
    assign c_out_15=g_0_15|(p_0_15&cin);
    assign c_out_16=g_0_16|(p_0_16&cin);
    assign c_out_17=g_0_17|(p_0_17&cin);
    assign c_out_18=g_0_18|(p_0_18&cin);
    assign c_out_19=g_0_19|(p_0_19&cin);
    assign c_out_20=g_0_20|(p_0_20&cin);
    assign c_out_21=g_0_21|(p_0_21&cin);
    assign c_out_22=g_0_22|(p_0_22&cin);
    assign c_out_23=g_0_23|(p_0_23&cin);
    assign c_out_24=g_0_24|(p_0_24&cin);
    assign c_out_25=g_0_25|(p_0_25&cin);
    assign c_out_26=g_0_26|(p_0_26&cin);
    assign c_out_27=g_0_27|(p_0_27&cin);
    assign c_out_28=g_0_28|(p_0_28&cin);
    assign c_out_29=g_0_29|(p_0_29&cin);
    assign c_out_30=g_0_30|(p_0_30&cin);
    assign c_out_31=g_0_31|(p_0_31&cin);
    assign sum[0]=p_0_0^cin;
    assign sum[1]=p_1_1^c_out_0;
    assign sum[2]=p_2_2^c_out_1;
    assign sum[3]=p_3_3^c_out_2;
    assign sum[4]=p_4_4^c_out_3;
    assign sum[5]=p_5_5^c_out_4;
    assign sum[6]=p_6_6^c_out_5;
    assign sum[7]=p_7_7^c_out_6;
    assign sum[8]=p_8_8^c_out_7;
    assign sum[9]=p_9_9^c_out_8;
    assign sum[10]=p_10_10^c_out_9;
    assign sum[11]=p_11_11^c_out_10;
    assign sum[12]=p_12_12^c_out_11;
    assign sum[13]=p_13_13^c_out_12;
    assign sum[14]=p_14_14^c_out_13;
    assign sum[15]=p_15_15^c_out_14;
    assign sum[16]=p_16_16^c_out_15;
    assign sum[17]=p_17_17^c_out_16;
    assign sum[18]=p_18_18^c_out_17;
    assign sum[19]=p_19_19^c_out_18;
    assign sum[20]=p_20_20^c_out_19;
    assign sum[21]=p_21_21^c_out_20;
    assign sum[22]=p_22_22^c_out_21;
    assign sum[23]=p_23_23^c_out_22;
    assign sum[24]=p_24_24^c_out_23;
    assign sum[25]=p_25_25^c_out_24;
    assign sum[26]=p_26_26^c_out_25;
    assign sum[27]=p_27_27^c_out_26;
    assign sum[28]=p_28_28^c_out_27;
    assign sum[29]=p_29_29^c_out_28;
    assign sum[30]=p_30_30^c_out_29;
    assign sum[31]=p_31_31^c_out_30;
    assign carryOut=c_out_31;
    assign overflow = c_out_31 ^ c_out_30;
    assign zero = (sum == 32'b0);
    assign neg = sum[31];
endmodule
